library verilog;
use verilog.vl_types.all;
entity Lab9_2_vlg_vec_tst is
end Lab9_2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Lab1_2_vlg_check_tst is
    port(
        carry           : in     vl_logic;
        S1              : in     vl_logic;
        S2              : in     vl_logic;
        S3              : in     vl_logic;
        S4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab1_2_vlg_check_tst;

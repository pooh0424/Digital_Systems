library verilog;
use verilog.vl_types.all;
entity Lab2_1_1_vlg_vec_tst is
end Lab2_1_1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Lab9_1_vlg_vec_tst is
end Lab9_1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Lab8_1_vlg_vec_tst is
end Lab8_1_vlg_vec_tst;

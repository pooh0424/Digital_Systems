library verilog;
use verilog.vl_types.all;
entity Lab6_1_vlg_sample_tst is
    port(
        KEY             : in     vl_logic_vector(2 downto 1);
        sampler_tx      : out    vl_logic
    );
end Lab6_1_vlg_sample_tst;

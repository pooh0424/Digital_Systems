library verilog;
use verilog.vl_types.all;
entity Lab3_1_vlg_check_tst is
    port(
        sevensegement   : in     vl_logic_vector(0 to 6);
        sampler_rx      : in     vl_logic
    );
end Lab3_1_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Lab12_1_vlg_vec_tst is
end Lab12_1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Lab8_2_vlg_vec_tst is
end Lab8_2_vlg_vec_tst;

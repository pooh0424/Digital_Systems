Library IEEE;
use IEEE.STD_Logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY Vbar_display IS   
	PORT( video_on:IN std_logic;
          r,c: IN INTEGER RANGE 0 TO 799;
		  Rout, Gout, Bout: out std_logic_vector(3 downto 0);
		  switch:IN std_logic_vector(5 downto 0));
END Vbar_display;

ARCHITECTURE arch OF Vbar_display IS
	constant circle:std_logic_vector(0 to 9799):=x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555575555555555555555555555555555555FFFFFFFD55555555555555555555555557FFFFFFFFFF55555555555555555555555FFFFFFFFFFFFFD555555555555555555557FFFFFFFFFFFFFF55555555555555555557FFFFFFFFFFFFFFFF555555555555555557FFFFFFFFFFFFFFFFFF5555555555555555FFFFFFFFFFFFFFFFFFFD555555555555557FFFFFFFFFFFFFFFFFFFF55555555555555FFFFFFFFFFFFFFFFFFFFFD5555555555557FFFFFFFFFFFFFFFFFFFFFF555555555555FFFFFFFFFFFFFFFFFFFFFFFD55555555557FFFFFFFFFFFFFFFFFFFFFFFF55555555557FFFFFFFFFFFFFFFFFFFFFFFF5555555555FFFFFFFFFFFFFFFFFFFFFFFFFD555555555FFFFFFFFFFFFFFFFFFFFFFFFFD555555557FFFFFFFFFFFFFFFFFFFFFFFFFF55555555FFFFFFFFFFFFFFFFFFFFFFFFFFFD5555555FFFFFFFFFFFFFFFFFFFFFFFFFFFD5555555FFFFFFFFFFFFFFFFFFFFFFFFFFFD5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFF5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFF5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFF555555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555557FFFFFFFFFFFFFFFFFFFFFFFFFFFF5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFF5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFF5555555FFFFFFFFFFFFFFFFFFFFFFFFFFFD5555555FFFFFFFFFFFFFFFFFFFFFFFFFFFD5555555FFFFFFFFFFFFFFFFFFFFFFFFFFFD55555557FFFFFFFFFFFFFFFFFFFFFFFFFF555555555FFFFFFFFFFFFFFFFFFFFFFFFFD555555555FFFFFFFFFFFFFFFFFFFFFFFFFD5555555557FFFFFFFFFFFFFFFFFFFFFFFF55555555557FFFFFFFFFFFFFFFFFFFFFFFF55555555555FFFFFFFFFFFFFFFFFFFFFFFD555555555557FFFFFFFFFFFFFFFFFFFFFF5555555555555FFFFFFFFFFFFFFFFFFFFFD55555555555557FFFFFFFFFFFFFFFFFFFF555555555555555FFFFFFFFFFFFFFFFFFFD5555555555555557FFFFFFFFFFFFFFFFFF555555555555555557FFFFFFFFFFFFFFFF55555555555555555557FFFFFFFFFFFFFF555555555555555555555FFFFFFFFFFFFFD55555555555555555555557FFFFFFFFFF55555555555555555555555555FFFFFFFD55555555555555555555555555555575555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555";

	constant le:std_logic_vector(0 to 9799):=x"555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555565555555555555555555555555555555AAAAAAA955555555555555555555555556AAAAAAAAAA55555555555555555555555AAAAAAAAAAAAA9555555555555555555556AAAAAAAAAAAAAA55555555555555555556AAAAAAAAAAAAAAAA555555555555555556AAAAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAAAAA9555555555555556AAAAAAAAAAAAAAAAAAAA55555555555555AAAAAAAAAAAAAAAAAAAAA95555555555556AAAAAAAAAABAAAAAAAAAAA555555555555AAAAAAAAAAAFEAAAAAAAAAA955555555556AAAAAAAAAABFFAAAAAAAAAAA55555555556AAAAAAAAAAFFEAAAAAAAAAAA5555555555AAAAAAAAAABFFAAAAAAAAAAAA9555555555AAAAAAAAAAFFEAAAAAAAAAAAA9555555556AAAAAAAAABFFAAAAAAAAAAAAAA55555555AAAAAAAAAAFFEAAAAAAAAAAAAAA95555555AAAAAAAAABFFAAAAAAAAAAAAAAA95555555AAAAAAAAAFFEAAAAAAAAAAAAAAA95555556AAAAAAAABFFAAAAAAAAAAAAAAAAA5555556AAAAAAAAFFEAAAAAAAAAAAAAAAAA5555556AAAAAAABFFAAAAAAAAAAAAAAAAAA555555AAAAAAAAFFEAAAAAAAAAAAAAAAAAA955555AAAAAAABFFAAAAAAAAAAAAAAAAAAA955555AAAAAAAFFEAAAAAAAAAAAAAAAAAAA955555AAAAAABFFAAAAAAAAAAAAAAAAAAAA955555AAAAAAFFEAAAAAAAAAAAAAAAAAAAA955555AAAAABFFAAAAAAAAAAAAAAAAAAAAA955555AAAAAFFEAAABFFFFFFFFFFFFAAAAA955556AAAABFFAAAABFFFFFFFFFFFFAAAAAA55555AAAAAFFEAAABFFFFFFFFFFFFAAAAA955555AAAAABFFAAABFFFFFFFFFFFFAAAAA955555AAAAAAFFEAAAAAAAAAAAAAAAAAAAA955555AAAAAABFFAAAAAAAAAAAAAAAAAAAA955555AAAAAAAFFEAAAAAAAAAAAAAAAAAAA955555AAAAAAABFFAAAAAAAAAAAAAAAAAAA955555AAAAAAAAFFEAAAAAAAAAAAAAAAAAA9555556AAAAAAABFFAAAAAAAAAAAAAAAAAA5555556AAAAAAAAFFEAAAAAAAAAAAAAAAAA5555556AAAAAAAABFFAAAAAAAAAAAAAAAAA5555555AAAAAAAAAFFEAAAAAAAAAAAAAAA95555555AAAAAAAAABFFAAAAAAAAAAAAAAA95555555AAAAAAAAAAFFEAAAAAAAAAAAAAA955555556AAAAAAAAABFFAAAAAAAAAAAAAA555555555AAAAAAAAAAFFEAAAAAAAAAAAA9555555555AAAAAAAAAABFFAAAAAAAAAAAA95555555556AAAAAAAAAAFFEAAAAAAAAAAA55555555556AAAAAAAAAABFFAAAAAAAAAAA55555555555AAAAAAAAAAAFEAAAAAAAAAA9555555555556AAAAAAAAAABAAAAAAAAAAA5555555555555AAAAAAAAAAAAAAAAAAAAA955555555555556AAAAAAAAAAAAAAAAAAAA555555555555555AAAAAAAAAAAAAAAAAAA95555555555555556AAAAAAAAAAAAAAAAAA555555555555555556AAAAAAAAAAAAAAAA55555555555555555556AAAAAAAAAAAAAA555555555555555555555AAAAAAAAAAAAA955555555555555555555556AAAAAAAAAA55555555555555555555555555AAAAAAA95555555555555555555555555555556555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555";
	constant ce:std_logic_vector(0 to 9799):=x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555565555555555555555555555555555555AAAAAAA955555555555555555555555556AAAAAAAAAA55555555555555555555555AAAAAAAAAAAAA9555555555555555555556AAAAAAAAAAAAAA55555555555555555556AAAAAAAAAAAAAAAA555555555555555556AAAAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAAAAA9555555555555556AAAAAAAAAAAAAAAAAAAA55555555555555AAAAAAAAAAAAAAAAAAAAA95555555555556AAAAAAAAAABAAAAAAAAAAA555555555555AAAAAAAAAAAFEAAAAAAAAAA955555555556AAAAAAAAAABFFAAAAAAAAAAA55555555556AAAAAAAAAAFFFEAAAAAAAAAA5555555555AAAAAAAAAABFFFFAAAAAAAAAA9555555555AAAAAAAAAAFFEFFEAAAAAAAAA9555555556AAAAAAAAABFFABFFAAAAAAAAAA55555555AAAAAAAAAAFFEAAFFEAAAAAAAAA95555555AAAAAAAAABFFAAABFFAAAAAAAAA95555555AAAAAAAAAFFEAAAAFFEAAAAAAAA95555556AAAAAAAABFFAAAAABFFAAAAAAAAA5555556AAAAAAAAFFEAAAAAAFFEAAAAAAAA5555556AAAAAAABFFAAAAAAABFFAAAAAAAA555555AAAAAAAAFFEAAAAAAAAFFEAAAAAAA955555AAAAAAABFFAAABFEAAABFFAAAAAAA955555AAAAAAAFFEAAABFEAAAAFFEAAAAAA955555AAAAAABFFAAAABFEAAAABFFAAAAAA955555AAAAAAFFEAAAABFEAAAAAFFEAAAAA955555AAAAABFFAAAAABFEAAAAABFFAAAAA955555AAAAAFFEAAAAABFEAAAAAAFFEAAAA955556AAAABFFAAAAAABFEAAAAAABFFAAAAA55555AAAAAFEAAAAAABFEAAAAAAAFEAAAA955555AAAAABAAAAAAABFEAAAAAAABAAAAA955555AAAAAAAAAAAAABFEAAAAAAAAAAAAA955555AAAAAAAAAAAAABFEAAAAAAAAAAAAA955555AAAAAAAAAAAAABFEAAAAAAAAAAAAA955555AAAAAAAAAAAAABFEAAAAAAAAAAAAA955555AAAAAAAAAAAAABFEAAAAAAAAAAAAA9555556AAAAAAAAAAAABFEAAAAAAAAAAAAA5555556AAAAAAAAAAAABFEAAAAAAAAAAAAA5555556AAAAAAAAAAAABFEAAAAAAAAAAAAA5555555AAAAAAAAAAAABFEAAAAAAAAAAAA95555555AAAAAAAAAAAABFEAAAAAAAAAAAA95555555AAAAAAAAAAAABFEAAAAAAAAAAAA955555556AAAAAAAAAAABFEAAAAAAAAAAAA555555555AAAAAAAAAAABFEAAAAAAAAAAA9555555555AAAAAAAAAAABFEAAAAAAAAAAA95555555556AAAAAAAAAABFEAAAAAAAAAAA55555555556AAAAAAAAAABFEAAAAAAAAAAA55555555555AAAAAAAAAAAAAAAAAAAAAAA9555555555556AAAAAAAAAAAAAAAAAAAAAA5555555555555AAAAAAAAAAAAAAAAAAAAA955555555555556AAAAAAAAAAAAAAAAAAAA555555555555555AAAAAAAAAAAAAAAAAAA95555555555555556AAAAAAAAAAAAAAAAAA555555555555555556AAAAAAAAAAAAAAAA55555555555555555556AAAAAAAAAAAAAA555555555555555555555AAAAAAAAAAAAA955555555555555555555556AAAAAAAAAA55555555555555555555555555AAAAAAA955555555555555555555555555555565555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555";
	constant ri:std_logic_vector(0 to 9799):=x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555595555555555555555555555555555556AAAAAAA55555555555555555555555555AAAAAAAAAA955555555555555555555556AAAAAAAAAAAAA555555555555555555555AAAAAAAAAAAAAA95555555555555555555AAAAAAAAAAAAAAAA955555555555555555AAAAAAAAAAAAAAAAAA95555555555555556AAAAAAAAAAAAAAAAAAA555555555555555AAAAAAAAAAAAAAAAAAAA955555555555556AAAAAAAAAAAAAAAAAAAAA5555555555555AAAAAAAAAAAEAAAAAAAAAA9555555555556AAAAAAAAAABFAAAAAAAAAAA55555555555AAAAAAAAAAAFFEAAAAAAAAAA95555555555AAAAAAAAAAABFFAAAAAAAAAA95555555556AAAAAAAAAAAAFFEAAAAAAAAAA5555555556AAAAAAAAAAAABFFAAAAAAAAAA555555555AAAAAAAAAAAAAAFFEAAAAAAAAA955555556AAAAAAAAAAAAAABFFAAAAAAAAAA55555556AAAAAAAAAAAAAAAFFEAAAAAAAAA55555556AAAAAAAAAAAAAAABFFAAAAAAAAA5555555AAAAAAAAAAAAAAAAAFFEAAAAAAAA9555555AAAAAAAAAAAAAAAAABFFAAAAAAAA9555555AAAAAAAAAAAAAAAAAAFFEAAAAAAA9555556AAAAAAAAAAAAAAAAAABFFAAAAAAAA555556AAAAAAAAAAAAAAAAAAAFFEAAAAAAA555556AAAAAAAAAAAAAAAAAAABFFAAAAAAA555556AAAAAAAAAAAAAAAAAAAAFFEAAAAAA555556AAAAAAAAAAAAAAAAAAAABFFAAAAAA555556AAAAAFFFFFFFFFFFFEAAAFFEAAAAA555556AAAAAFFFFFFFFFFFFEAAABFFAAAAA55555AAAAAAFFFFFFFFFFFFEAAAAFFEAAAA955556AAAAAFFFFFFFFFFFFEAAABFFAAAAA555556AAAAAAAAAAAAAAAAAAAAAFFEAAAAA555556AAAAAAAAAAAAAAAAAAAABFFAAAAAA555556AAAAAAAAAAAAAAAAAAAAFFEAAAAAA555556AAAAAAAAAAAAAAAAAAABFFAAAAAAA555556AAAAAAAAAAAAAAAAAAAFFEAAAAAAA555556AAAAAAAAAAAAAAAAAABFFAAAAAAAA555555AAAAAAAAAAAAAAAAAAFFEAAAAAAA9555555AAAAAAAAAAAAAAAAABFFAAAAAAAA9555555AAAAAAAAAAAAAAAAAFFEAAAAAAAA95555556AAAAAAAAAAAAAAABFFAAAAAAAAA55555556AAAAAAAAAAAAAAAFFEAAAAAAAAA55555556AAAAAAAAAAAAAABFFAAAAAAAAAA55555555AAAAAAAAAAAAAAFFEAAAAAAAAA9555555556AAAAAAAAAAAABFFAAAAAAAAAA5555555556AAAAAAAAAAAAFFEAAAAAAAAAA5555555555AAAAAAAAAAABFFAAAAAAAAAA95555555555AAAAAAAAAAAFFEAAAAAAAAAA955555555556AAAAAAAAAABFAAAAAAAAAAA555555555555AAAAAAAAAAAEAAAAAAAAAA95555555555556AAAAAAAAAAAAAAAAAAAAA55555555555555AAAAAAAAAAAAAAAAAAAA9555555555555556AAAAAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAAAA955555555555555555AAAAAAAAAAAAAAAA95555555555555555555AAAAAAAAAAAAAA9555555555555555555556AAAAAAAAAAAAA55555555555555555555555AAAAAAAAAA955555555555555555555555556AAAAAAA555555555555555555555555555555595555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555";
begin
process(video_on,r,c) 
variable nowpos:IntEGER;
begin
If video_on='1' then         
    IF (r>=0 AND r<210)and (c>=0 and c<210) THEN
		nowpos:=(r/3*70+c/3)*2;
	   if circle(nowpos to nowpos+1)="01" then
			Rout<="1111"; Gout<="1111"; Bout<="1111";
		elsif circle(nowpos to nowpos+1)="10" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		elsif circle(nowpos to nowpos+1)="11"and switch(5)='1' then
			Rout<="1111"; Gout<="0000"; Bout<="0000";
		elsif circle(nowpos to nowpos+1)="11" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		end if;
	 elsif (r>=0 AND r<210) and (c>=210 and c<420) THEN
		nowpos:=(r/3*70+(c-210)/3)*2;
	   if circle(nowpos to nowpos+1)="01" then
			Rout<="1111"; Gout<="1111"; Bout<="1111";
		elsif circle(nowpos to nowpos+1)="10" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		elsif circle(nowpos to nowpos+1)="11" and switch(4)='1' then
			Rout<="1111"; Gout<="1111"; Bout<="0000";
		elsif circle(nowpos to nowpos+1)="11" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		end if;
	 elsif (r>=0 AND r<210) and (c>=420 and c<630)  THEN
		nowpos:=(r/3*70+(c-420)/3)*2;
	   if circle(nowpos to nowpos+1)="01" then
			Rout<="1111"; Gout<="1111"; Bout<="1111";
		elsif circle(nowpos to nowpos+1)="10" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		elsif circle(nowpos to nowpos+1)="11"and switch(3)='1' then
			Rout<="0000"; Gout<="1111"; Bout<="0000";
		elsif circle(nowpos to nowpos+1)="11" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		end if;
    elsif (r>=210 AND r<420)and (c>=0 and c<210) THEN
		nowpos:=((r-210)/3*70+c/3)*2;
	   if le(nowpos to nowpos+1)="01" then
			Rout<="1111"; Gout<="1111"; Bout<="1111";
		elsif le(nowpos to nowpos+1)="10" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		elsif le(nowpos to nowpos+1)="11"and switch(2)='1' then
			Rout<="0000"; Gout<="1111"; Bout<="0000";
		elsif le(nowpos to nowpos+1)="11" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		end if;
	 elsif (r>=210 AND r<420) and (c>=210 and c<420) THEN
		nowpos:=((r-210)/3*70+(c-210)/3)*2;
	   if ce(nowpos to nowpos+1)="01" then
			Rout<="1111"; Gout<="1111"; Bout<="1111";
		elsif ce(nowpos to nowpos+1)="10" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		elsif ce(nowpos to nowpos+1)="11"and switch(1)='1' then
			Rout<="0000"; Gout<="1111"; Bout<="0000";
		elsif ce(nowpos to nowpos+1)="11" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		end if;
	 elsif (r>=210 AND r<420) and (c>=420 and c<630)  THEN
		nowpos:=((r-210)/3*70+(c-420)/3)*2;
	   if ri(nowpos to nowpos+1)="01" then
			Rout<="1111"; Gout<="1111"; Bout<="1111";
		elsif ri(nowpos to nowpos+1)="10" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		elsif ri(nowpos to nowpos+1)="11"and switch(0)='1' then
			Rout<="0000"; Gout<="1111"; Bout<="0000";
		elsif ri(nowpos to nowpos+1)="11" then
			Rout<="0000"; Gout<="0000"; Bout<="0000";
		end if;
    else
       Rout<="0000"; Gout<="0000"; Bout<="0000";
    end if;
	 
else                            
    Rout<="0000"; Gout<="0000"; Bout<="0000";
end if;
end process;

END arch;

library ieee;
use ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all ;
entity Lab4_2 is
	port (
		SW: in std_logic_vector(5 downto 0);
		KEY: in std_logic_vector(1 downto 0);
		HEX0: out std_logic_vector(0 to 6);
		HEX1: out std_logic_vector(0 to 6);
		LEDG: out std_logic_vector(3 downto 0)
	);
end  Lab4_2;
architecture behavor of Lab4_2 is
	SIGNAL SWA:std_logic_vector(3 downto 0);
	SIGNAL SWB:std_logic_vector(3 downto 0);
	SIGNAL SUM:std_logic_vector(3 downto 0);
begin
	SWA(2 downto 0)<=SW(5 downto 3);
	SWB(2 downto 0)<=SW(2 downto 0);
	PROCESS(KEY)
	BEGIN
		SUM<=SWA+SWB;
		IF KEY="10" THEN
			CASE SUM IS
				WHEN "0001" =>HEX0<="1001111" ;HEX1<="0000001";
				WHEN "0010" =>HEX0<="0010010" ;HEX1<="0000001";
				WHEN "0011" =>HEX0<="0000110" ;HEX1<="0000001";
				WHEN "0100" =>HEX0<="1001100" ;HEX1<="0000001";
				WHEN "0101" =>HEX0<="0100100" ;HEX1<="0000001";
				WHEN "0110" =>HEX0<="0100000" ;HEX1<="0000001";
				WHEN "0111" =>HEX0<="0001111" ;HEX1<="0000001";
				WHEN "1000" =>HEX0<="0000000" ;HEX1<="0000001";
				WHEN "1001" =>HEX0<="0001100" ;HEX1<="0000001";
				WHEN "1010" =>HEX0<="0000001" ;HEX1<="1001111";
				WHEN "1011" =>HEX0<="1001111" ;HEX1<="1001111";
				WHEN "1100" =>HEX0<="0010010" ;HEX1<="1001111";
				WHEN "1101" =>HEX0<="0000110" ;HEX1<="1001111";
				WHEN "1110" =>HEX0<="1001100" ;HEX1<="1001111";
				WHEN "1111" =>HEX0<="0100100" ;HEX1<="1001111";
				WHEN OTHERS =>HEX0<="0000001" ;HEX1<="0000001";
			END CASE;
		ELSIF KEY="01" THEN
			LEDG <= SUM;
		ELSE
			LEDG <= "0000";
			HEX0<="1111111";
			HEX1<="1111111";
		END IF;
	END PROCESS;
	
end behavor ;  

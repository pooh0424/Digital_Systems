library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
entity paritice3 is 
port(	CLOCK_50:in std_logic;
		SW:in std_LOGIC_Vector(5 downto 0);
		VGA_R, VGA_G, VGA_B: out std_logic_vector(3 downto 0);
		VGA_HS,VGA_VS: OUT std_logic
		);
end paritice3;

architecture behavor of paritice3 is
component VGA_sync IS
	PORT(
		CLOCK,RESET: IN std_logic;
		HOR_SYN,VER_SYN,video_on: OUT std_logic;
      row_counter:out INTEGER RANGE 0 TO 524;		
      col_counter:out INTEGER RANGE 0 TO 799	);
END component;
component Vbar_display IS   
	PORT( video_on:IN std_logic;
   r,c: IN INTEGER RANGE 0 TO 799;
	Rout, Gout, Bout: out std_logic_vector(3 downto 0);
	switch:in std_LOGIC_Vector(5 downto 0));
END component;

component CLK_DIV is
	port 
	(	
		clock_in				: IN	STD_LOGIC;
		clock_out			: OUT	STD_LOGIC); 
end component;
signal clock25:std_logic;
signal r,c:INTEGER RANGE 0 TO 799;
signal video_on:std_LOGIC;
begin
	VGA_sync1:VGA_sync port map(clock25,'1',VGA_HS,VGA_VS,video_on,r,c);
	Vbar_display1:Vbar_display port map(video_on,r,c,VGA_R,VGA_G,VGA_B,sw);
	clock_div1:CLK_DIV port map(cloCK_50,clock25);
end Behavor;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity CLK_DIV is
	port 
	(	
		clock_in				: IN	STD_LOGIC;
		clock_out			: OUT	STD_LOGIC); 
end CLK_DIV;

architecture arch of CLK_DIV is
	signal CLK_out: STD_LOGIC;
begin
	process(clock_in)
	begin
		IF clock_in'event and clock_in='1' THEN
				CLK_out <= NOT CLK_out;
		END IF;
		clock_out <= CLK_out;
	end process;
end arch;




library verilog;
use verilog.vl_types.all;
entity Lab1_2 is
    port(
        S1              : out    vl_logic;
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        M               : in     vl_logic;
        S2              : out    vl_logic;
        A2              : in     vl_logic;
        B2              : in     vl_logic;
        S3              : out    vl_logic;
        A3              : in     vl_logic;
        B3              : in     vl_logic;
        S4              : out    vl_logic;
        A4              : in     vl_logic;
        B4              : in     vl_logic;
        carry           : out    vl_logic
    );
end Lab1_2;
